module fft();

endmodule
