module randomizer(
	input reset, clk
	input in_bits,
	input in_valid,
	output out_bits,
	output out_valid
	input [14:0] rand_iv,
	input reload);

endmodule
