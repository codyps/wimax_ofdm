module cp(
	input reset, clk,
	input [1:0] param_G,
	input cp_in_bits,
	input cp_in_valid,
	output cp_out_bits,
	output cp_out_valid
	/* FIXME: these widths are probably wrong. */
);

endmodule
